* C:\Users\PREM\eSim-Workspace\notgatev1\notgatev1.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 02/10/22 00:54:10

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M2  /not_output /not_input GND GND mosfet_n		
M1  /not_output /not_input /vdd /vdd mosfet_p		
U1  /vdd /not_input /not_output PORT		

.end

* C:\Users\PREM\eSim-Workspace\andgatev1\andgatev1.cir
.lib "sky130_fd_pr/models/sky130.lib.spice" tt

*3 input AND
xM1  Net-_M1-Pad1_ in1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		
xM2  Net-_M1-Pad1_ in2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		
xM3  Net-_M1-Pad1_ ena vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		
xM4  Net-_M1-Pad1_ in1 Net-_M4-Pad3_ Net-_M4-Pad3_ sky130_fd_pr__nfet_01v8 w=.42 l=.5		
xM5  Net-_M4-Pad3_ in2 Net-_M5-Pad3_ Net-_M5-Pad3_ sky130_fd_pr__nfet_01v8 w=.42 l=.5		
xM6  Net-_M5-Pad3_ ena GND GND sky130_fd_pr__nfet_01v8 w=.42 l=.5		

*inverter		
xM8  out Net-_M1-Pad1_ GND GND sky130_fd_pr__nfet_01v8 w=.42 l=.5		
xM7  out Net-_M1-Pad1_ vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		

Vdd vdd 0 3.3
Vin_1 ena 0 3
Vd0 in1 0 pulse(0 3 0s 0s 0s 5us 10us)
Vd1 in2 0 pulse(0 3 0s 0s 0s 10us 20us)

.tran 0.1us 20us

.control
run
plot V(in1) V(in2)+5 V(out)+10 V(ena)+15
.endc
.end
